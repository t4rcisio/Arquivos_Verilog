






module clcok_manager(clock, clock_00, clock_01, clock_02, clock_03);