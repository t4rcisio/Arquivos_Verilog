library verilog;
use verilog.vl_types.all;
entity nRisc_core is
    port(
        clock           : in     vl_logic
    );
end nRisc_core;
